** Profile: "SCHEMATIC1-tf_pid_ramp"  [ C:\Program Files\Orcad\Files\tf_pid_ramp-SCHEMATIC1-tf_pid_ramp.sim ] 

** Creating circuit file "tf_pid_ramp-SCHEMATIC1-tf_pid_ramp.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tf_pid_ramp-SCHEMATIC1.net" 


.END
