** Profile: "SCHEMATIC1-DEL_recent"  [ C:\Program Files\Orcad\Files\del_recent-SCHEMATIC1-DEL_recent.sim ] 

** Creating circuit file "del_recent-SCHEMATIC1-DEL_recent.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\del_recent-SCHEMATIC1.net" 


.END
