** Profile: "SCHEMATIC1-parabola"  [ C:\Program Files\Orcad\Files\tf_pid_parab-SCHEMATIC1-parabola.sim ] 

** Creating circuit file "tf_pid_parab-SCHEMATIC1-parabola.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10s 0 SKIPBP 
.OPTIONS STEPGMIN
.OPTIONS ABSTOL= 1.0n
.OPTIONS ITL4= 100
.OPTIONS RELTOL= 0.01
.OPTIONS VNTOL= 1.0m
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tf_pid_parab-SCHEMATIC1.net" 


.END
