** Profile: "SCHEMATIC1-TF_RAMP"  [ C:\Program Files\Orcad\Files\tf_ramp-SCHEMATIC1-TF_RAMP.sim ] 

** Creating circuit file "tf_ramp-SCHEMATIC1-TF_RAMP.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 1.5 SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tf_ramp-SCHEMATIC1.net" 


.END
