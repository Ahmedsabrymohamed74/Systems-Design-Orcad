** Profile: "SCHEMATIC1-tf_parab"  [ C:\Program Files\Orcad\Files\tf_lag_parabolic_tune-SCHEMATIC1-tf_parab.sim ] 

** Creating circuit file "tf_lag_parabolic_tune-SCHEMATIC1-tf_parab.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 100k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tf_lag_parabolic_tune-SCHEMATIC1.net" 


.END
