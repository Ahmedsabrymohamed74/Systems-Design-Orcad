** Profile: "SCHEMATIC1-step_g"  [ C:\Program Files\Orcad\Files\g(s) -SCHEMATIC1-step_g.sim ] 

** Creating circuit file "g(s) -SCHEMATIC1-step_g.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000s 0 SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\g(s) -SCHEMATIC1.net" 


.END
