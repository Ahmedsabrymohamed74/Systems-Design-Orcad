** Profile: "SCHEMATIC1-parab_tfPid"  [ C:\Program Files\Orcad\Files\tf_pid_parab-SCHEMATIC1-parab_tfPid.sim ] 

** Creating circuit file "tf_pid_parab-SCHEMATIC1-parab_tfPid.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tf_pid_parab-SCHEMATIC1.net" 


.END
