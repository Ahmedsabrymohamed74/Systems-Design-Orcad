** Profile: "SCHEMATIC1-stepimp"  [ C:\Program Files\Orcad\Files\g(s)_impulse-SCHEMATIC1-stepimp.sim ] 

** Creating circuit file "g(s)_impulse-SCHEMATIC1-stepimp.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10s 0 SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\g(s)_impulse-SCHEMATIC1.net" 


.END
