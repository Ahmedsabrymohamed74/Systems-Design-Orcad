** Profile: "SCHEMATIC1-design1"  [ C:\Program Files\Orcad\Files\lag_designs-SCHEMATIC1-design1.sim ] 

** Creating circuit file "lag_designs-SCHEMATIC1-design1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lag_designs-SCHEMATIC1.net" 


.END
