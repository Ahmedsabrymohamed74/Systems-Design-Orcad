** Profile: "SCHEMATIC1-stepg"  [ C:\Program Files\Orcad\Files\g(s)_step-SCHEMATIC1-stepg.sim ] 

** Creating circuit file "g(s)_step-SCHEMATIC1-stepg.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10 0 SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\g(s)_step-SCHEMATIC1.net" 


.END
