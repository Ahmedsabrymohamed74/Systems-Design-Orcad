** Profile: "SCHEMATIC1-pidstep"  [ C:\Program Files\Orcad\Files\tf_pid_step-SCHEMATIC1-pidstep.sim ] 

** Creating circuit file "tf_pid_step-SCHEMATIC1-pidstep.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tf_pid_step-SCHEMATIC1.net" 


.END
